10'b100111_0100
10'b110101_0100
10'b100111_1001
10'b110101_1001
10'b100111_0101
10'b110101_0101
10'b100111_0011
10'b110101_0011
10'b100111_0010
10'b110101_0010
10'b100111_1010
10'b110101_1010
10'b100111_0110
10'b110101_0110
10'b100111_0001
10'b110101_0001
10'b011101_0100
10'b101001_1011
10'b011101_1001
10'b101001_1001
10'b011101_0101
10'b101001_0101
10'b011101_0011
10'b101001_1100
10'b011101_0010
10'b101001_1101
10'b011101_1010
10'b101001_1010
10'b011101_0110
10'b101001_0110
10'b011101_0001
10'b101001_1110
10'b101101_0100
10'b011001_1011
10'b101101_1001
10'b011001_1001
10'b101101_0101
10'b011001_0101
10'b101101_0011
10'b011001_1100
10'b101101_0010
10'b011001_1101
10'b101101_1010
10'b011001_1010
10'b101101_0110
10'b011001_0110
10'b101101_0001
10'b011001_1110
10'b110001_1011
10'b111000_1011
10'b110001_1001
10'b111000_1001
10'b110001_0101
10'b111000_0101
10'b110001_1100
10'b111000_1100
10'b110001_1101
10'b111000_1101
10'b110001_1010
10'b111000_1010
10'b110001_0110
10'b111000_0110
10'b110001_1110
10'b111000_1110
10'b111001_0100
10'b001101_1011
10'b111001_1001
10'b001101_1001
10'b111001_0101
10'b001101_0101
10'b111001_0011
10'b001101_1100
10'b111001_0010
10'b001101_1101
10'b111001_1010
10'b001101_1010
10'b111001_0110
10'b001101_0110
10'b111001_0001
10'b001101_1110
10'b100101_1011
10'b101100_1011
10'b100101_1001
10'b101100_1001
10'b100101_0101
10'b101100_0101
10'b100101_1100
10'b101100_1100
10'b100101_1101
10'b101100_1101
10'b100101_1010
10'b101100_1010
10'b100101_0110
10'b101100_0110
10'b100101_1110
10'b101100_1110
10'b010101_1011
10'b011100_1011
10'b010101_1001
10'b011100_1001
10'b010101_0101
10'b011100_0101
10'b010101_1100
10'b011100_1100
10'b010101_1101
10'b011100_1101
10'b010101_1010
10'b011100_1010
10'b010101_0110
10'b011100_0110
10'b010101_1110
10'b011100_1110
10'b110100_1011
10'b010111_0100
10'b110100_1001
10'b010111_1001
10'b110100_0101
10'b010111_0101
10'b110100_1100
10'b010111_0011
10'b110100_1101
10'b010111_0010
10'b110100_1010
10'b010111_1010
10'b110100_0110
10'b010111_0110
10'b110100_1110
10'b010111_0001
10'b011011_0100
10'b001011_1011
10'b011011_1001
10'b001011_1001
10'b011011_0101
10'b001011_0101
10'b011011_0011
10'b001011_1100
10'b011011_0010
10'b001011_1101
10'b011011_1010
10'b001011_1010
10'b011011_0110
10'b001011_0110
10'b011011_0001
10'b001011_0111
10'b100011_1011
10'b101010_1011
10'b100011_1001
10'b101010_1001
10'b100011_0101
10'b101010_0101
10'b100011_1100
10'b101010_1100
10'b100011_1101
10'b101010_1101
10'b100011_1010
10'b101010_1010
10'b100011_0110
10'b101010_0110
10'b100011_0111
10'b101010_1110
10'b010011_1011
10'b011010_1011
10'b010011_1001
10'b011010_1001
10'b010011_0101
10'b011010_0101
10'b010011_1100
10'b011010_1100
10'b010011_1101
10'b011010_1101
10'b010011_1010
10'b011010_1010
10'b010011_0110
10'b011010_0110
10'b010011_0111
10'b011010_1110
10'b110010_1011
10'b111010_0100
10'b110010_1001
10'b111010_1001
10'b110010_0101
10'b111010_0101
10'b110010_1100
10'b111010_0011
10'b110010_1101
10'b111010_0010
10'b110010_1010
10'b111010_1010
10'b110010_0110
10'b111010_0110
10'b110010_1110
10'b111010_0001
10'b110011_0100
10'b001110_1011
10'b110011_1001
10'b001110_1001
10'b110011_0101
10'b001110_0101
10'b110011_0011
10'b001110_1100
10'b110011_0010
10'b001110_1101
10'b110011_1010
10'b001110_1010
10'b110011_0110
10'b001110_0110
10'b110011_0001
10'b001110_1110
10'b100110_1011
10'b101110_0100
10'b100110_1001
10'b101110_1001
10'b100110_0101
10'b101110_0101
10'b100110_1100
10'b101110_0011
10'b100110_1101
10'b101110_0010
10'b100110_1010
10'b101110_1010
10'b100110_0110
10'b101110_0110
10'b100110_1110
10'b101110_0001
10'b010110_1011
10'b011110_0100
10'b010110_1001
10'b011110_1001
10'b010110_0101
10'b011110_0101
10'b010110_1100
10'b011110_0011
10'b010110_1101
10'b011110_0010
10'b010110_1010
10'b011110_1010
10'b010110_0110
10'b011110_0110
10'b010110_1110
10'b011110_0001
10'b110110_0100
10'b101011_0100
10'b110110_1001
10'b101011_1001
10'b110110_0101
10'b101011_0101
10'b110110_0011
10'b101011_0011
10'b110110_0010
10'b101011_0010
10'b110110_1010
10'b101011_1010
10'b110110_0110
10'b101011_0110
10'b110110_0001
10'b101011_0001
