10'b011000_1011
10'b001010_1011
10'b011000_1001
10'b001010_1001
10'b011000_0101
10'b001010_0101
10'b011000_1100
10'b001010_1100
10'b011000_1101
10'b001010_1101
10'b011000_1010
10'b001010_1010
10'b011000_0110
10'b001010_0110
10'b011000_1110
10'b001010_1110
10'b100010_1011
10'b101001_0100
10'b100010_1001
10'b101001_1001
10'b100010_0101
10'b101001_0101
10'b100010_1100
10'b101001_0011
10'b100010_1101
10'b101001_0010
10'b100010_1010
10'b101001_1010
10'b100010_0110
10'b101001_0110
10'b100010_1110
10'b101001_0001
10'b010010_1011
10'b011001_0100
10'b010010_1001
10'b011001_1001
10'b010010_0101
10'b011001_0101
10'b010010_1100
10'b011001_0011
10'b010010_1101
10'b011001_0010
10'b010010_1010
10'b011001_1010
10'b010010_0110
10'b011001_0110
10'b010010_1110
10'b011001_0001
10'b110001_0100
10'b000111_0100
10'b110001_1001
10'b000111_1001
10'b110001_0101
10'b000111_0101
10'b110001_0011
10'b000111_0011
10'b110001_0010
10'b000111_0010
10'b110001_1010
10'b000111_1010
10'b110001_0110
10'b000111_0110
10'b110001_0001
10'b000111_0001
10'b000110_1011
10'b001101_0100
10'b000110_1001
10'b001101_1001
10'b000110_0101
10'b001101_0101
10'b000110_1100
10'b001101_0011
10'b000110_1101
10'b001101_0010
10'b000110_1010
10'b001101_1010
10'b000110_0110
10'b001101_0110
10'b000110_1110
10'b001101_0001
10'b100101_0100
10'b101100_0100
10'b100101_1001
10'b101100_1001
10'b100101_0101
10'b101100_0101
10'b100101_0011
10'b101100_0011
10'b100101_0010
10'b101100_0010
10'b100101_1010
10'b101100_1010
10'b100101_0110
10'b101100_0110
10'b100101_0001
10'b101100_1000
10'b010101_0100
10'b011100_0100
10'b010101_1001
10'b011100_1001
10'b010101_0101
10'b011100_0101
10'b010101_0011
10'b011100_0011
10'b010101_0010
10'b011100_0010
10'b010101_1010
10'b011100_1010
10'b010101_0110
10'b011100_0110
10'b010101_0001
10'b011100_1000
10'b110100_0100
10'b101000_1011
10'b110100_1001
10'b101000_1001
10'b110100_0101
10'b101000_0101
10'b110100_0011
10'b101000_1100
10'b110100_0010
10'b101000_1101
10'b110100_1010
10'b101000_1010
10'b110100_0110
10'b101000_0110
10'b110100_1000
10'b101000_1110
10'b100100_1011
10'b001011_0100
10'b100100_1001
10'b001011_1001
10'b100100_0101
10'b001011_0101
10'b100100_1100
10'b001011_0011
10'b100100_1101
10'b001011_0010
10'b100100_1010
10'b001011_1010
10'b100100_0110
10'b001011_0110
10'b100100_1110
10'b001011_0001
10'b100011_0100
10'b101010_0100
10'b100011_1001
10'b101010_1001
10'b100011_0101
10'b101010_0101
10'b100011_0011
10'b101010_0011
10'b100011_0010
10'b101010_0010
10'b100011_1010
10'b101010_1010
10'b100011_0110
10'b101010_0110
10'b100011_0001
10'b101010_0001
10'b010011_0100
10'b011010_0100
10'b010011_1001
10'b011010_1001
10'b010011_0101
10'b011010_0101
10'b010011_0011
10'b011010_0011
10'b010011_0010
10'b011010_0010
10'b010011_1010
10'b011010_1010
10'b010011_0110
10'b011010_0110
10'b010011_0001
10'b011010_0001
10'b110010_0100
10'b000101_1011
10'b110010_1001
10'b000101_1001
10'b110010_0101
10'b000101_0101
10'b110010_0011
10'b000101_1100
10'b110010_0010
10'b000101_1101
10'b110010_1010
10'b000101_1010
10'b110010_0110
10'b000101_0110
10'b110010_0001
10'b000101_1110
10'b001100_1011
10'b001110_0100
10'b001100_1001
10'b001110_1001
10'b001100_0101
10'b001110_0101
10'b001100_1100
10'b001110_0011
10'b001100_1101
10'b001110_0010
10'b001100_1010
10'b001110_1010
10'b001100_0110
10'b001110_0110
10'b001100_1110
10'b001110_0001
10'b100110_0100
10'b010001_1011
10'b100110_1001
10'b010001_1001
10'b100110_0101
10'b010001_0101
10'b100110_0011
10'b010001_1100
10'b100110_0010
10'b010001_1101
10'b100110_1010
10'b010001_1010
10'b100110_0110
10'b010001_0110
10'b100110_0001
10'b010001_1110
10'b010110_0100
10'b100001_1011
10'b010110_1001
10'b100001_1001
10'b010110_0101
10'b100001_0101
10'b010110_0011
10'b100001_1100
10'b010110_0010
10'b100001_1101
10'b010110_1010
10'b100001_1010
10'b010110_0110
10'b100001_0110
10'b010110_0001
10'b100001_1110
10'b001001_1011
10'b010100_1011
10'b001001_1001
10'b010100_1001
10'b001001_0101
10'b010100_0101
10'b001001_1100
10'b010100_1100
10'b001001_1101
10'b010100_1101
10'b001001_1010
10'b010100_1010
10'b001001_0110
10'b010100_0110
10'b001001_1110
10'b010100_1110
