`include "crc32.v"
`include "enc3to4.v"
`include "enc5to6.v"
`include "kcode8to10.v"
`include "runningDisparity.v"
`include "enc8to10.v"


