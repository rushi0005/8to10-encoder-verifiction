class my_monitor_crc_in_message;

	logic pushin;
	logic [8:0] datain;
	logic startin;

endclass : my_monitor_crc_in_message
