class crc_output_packet;
	logic [39:0] crc_out;
endclass : crc_output_packet
