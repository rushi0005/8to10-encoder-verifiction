class my_monitor_crc_out_message;

	logic       pushout  ;//
	logic [9:0] dataout  ;//
	logic       startout ;
endclass : my_monitor_crc_out_message
