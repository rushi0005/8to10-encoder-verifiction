8'b000_00000
8'b000_00100
8'b001_00000
8'b001_00100
8'b010_00000
8'b010_00100
8'b011_00000
8'b011_00100
8'b100_00000
8'b100_00100
8'b101_00000
8'b101_00100
8'b110_00000
8'b110_00100
8'b111_00000
8'b111_00100
8'b000_00001
8'b000_00101
8'b001_00001
8'b001_00101
8'b010_00001
8'b010_00101
8'b011_00001
8'b011_00101
8'b100_00001
8'b100_00101
8'b101_00001
8'b101_00101
8'b110_00001
8'b110_00101
8'b111_00001
8'b111_00101
8'b000_00010
8'b000_00110
8'b001_00010
8'b001_00110
8'b010_00010
8'b010_00110
8'b011_00010
8'b011_00110
8'b100_00010
8'b100_00110
8'b101_00010
8'b101_00110
8'b110_00010
8'b110_00110
8'b111_00010
8'b111_00110
8'b000_00011
8'b000_00111
8'b001_00011
8'b001_00111
8'b010_00011
8'b010_00111
8'b011_00011
8'b011_00111
8'b100_00011
8'b100_00111
8'b101_00011
8'b101_00111
8'b110_00011
8'b110_00111
8'b111_00011
8'b111_00111
8'b000_01000
8'b000_01100
8'b001_01000
8'b001_01100
8'b010_01000
8'b010_01100
8'b011_01000
8'b011_01100
8'b100_01000
8'b100_01100
8'b101_01000
8'b101_01100
8'b110_01000
8'b110_01100
8'b111_01000
8'b111_01100
8'b000_01001
8'b000_01101
8'b001_01001
8'b001_01101
8'b010_01001
8'b010_01101
8'b011_01001
8'b011_01101
8'b100_01001
8'b100_01101
8'b101_01001
8'b101_01101
8'b110_01001
8'b110_01101
8'b111_01001
8'b111_01101
8'b000_01010
8'b000_01110
8'b001_01010
8'b001_01110
8'b010_01010
8'b010_01110
8'b011_01010
8'b011_01110
8'b100_01010
8'b100_01110
8'b101_01010
8'b101_01110
8'b110_01010
8'b110_01110
8'b111_01010
8'b111_01110
8'b000_01011
8'b000_01111
8'b001_01011
8'b001_01111
8'b010_01011
8'b010_01111
8'b011_01011
8'b011_01111
8'b100_01011
8'b100_01111
8'b101_01011
8'b101_01111
8'b110_01011
8'b110_01111
8'b111_01011
8'b111_01111
8'b000_10000
8'b000_10100
8'b001_10000
8'b001_10100
8'b010_10000
8'b010_10100
8'b011_10000
8'b011_10100
8'b100_10000
8'b100_10100
8'b101_10000
8'b101_10100
8'b110_10000
8'b110_10100
8'b111_10000
8'b111_10100
8'b000_10001
8'b000_10101
8'b001_10001
8'b001_10101
8'b010_10001
8'b010_10101
8'b011_10001
8'b011_10101
8'b100_10001
8'b100_10101
8'b101_10001
8'b101_10101
8'b110_10001
8'b110_10101
8'b111_10001
8'b111_10101
8'b000_10010
8'b000_10110
8'b001_10010
8'b001_10110
8'b010_10010
8'b010_10110
8'b011_10010
8'b011_10110
8'b100_10010
8'b100_10110
8'b101_10010
8'b101_10110
8'b110_10010
8'b110_10110
8'b111_10010
8'b111_10110
8'b000_10011
8'b000_10111
8'b001_10011
8'b001_10111
8'b010_10011
8'b010_10111
8'b011_10011
8'b011_10111
8'b100_10011
8'b100_10111
8'b101_10011
8'b101_10111
8'b110_10011
8'b110_10111
8'b111_10011
8'b111_10111
8'b000_11000
8'b000_11100
8'b001_11000
8'b001_11100
8'b010_11000
8'b010_11100
8'b011_11000
8'b011_11100
8'b100_11000
8'b100_11100
8'b101_11000
8'b101_11100
8'b110_11000
8'b110_11100
8'b111_11000
8'b111_11100
8'b000_11001
8'b000_11101
8'b001_11001
8'b001_11101
8'b010_11001
8'b010_11101
8'b011_11001
8'b011_11101
8'b100_11001
8'b100_11101
8'b101_11001
8'b101_11101
8'b110_11001
8'b110_11101
8'b111_11001
8'b111_11101
8'b000_11010
8'b000_11110
8'b001_11010
8'b001_11110
8'b010_11010
8'b010_11110
8'b011_11010
8'b011_11110
8'b100_11010
8'b100_11110
8'b101_11010
8'b101_11110
8'b110_11010
8'b110_11110
8'b111_11010
8'b111_11110
8'b000_11011
8'b000_11111
8'b001_11011
8'b001_11111
8'b010_11011
8'b010_11111
8'b011_11011
8'b011_11111
8'b100_11011
8'b100_11111
8'b101_11011
8'b101_11111
8'b110_11011
8'b110_11111
8'b111_11011
8'b111_11111


00011100001111_0100110000_1011
00111100001111_1001110000_0110
01011100001111_0101110000_1010
01111100001111_0011110000_1100
10011100001111_0010110000_1101
10111100001111_1010110000_0101
11011100001111_0110110000_1001
11111100001111_1000110000_0111
11110111111010_1000000101_0111
11111011110110_1000001001_0111
11111101101110_1000010001_0111
11111110011110_1000100001_0111
